// Verilog file written by procedure Aig_ManDumpVerilog()
module test ( n01, n02, n03, n04, n05, n06, n07, n08, n09, n10, n11, n12, n13, n14, n15, n16, n17 );
input n01;
input n02;
input n03;
input n04;
input n05;
input n06;
input n07;
input n08;
input n09;
input n10;
input n11;
input n12;
input n13;
input n14;
input n15;
input n16;
output n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
assign n18 =  n02 &  n04;
assign n19 = ~n07 & ~n10;
assign n20 = ~n05 & ~n09;
assign n21 = ~n19 & ~n20;
assign n22 = ~n11 & ~n21;
assign n23 = ~n06 & ~n08;
assign n24 = ~n22 &  n23;
assign n25 = ~n18 & ~n24;
assign n26 =  n08 &  n09;
assign n27 =  n05 & ~n08;
assign n28 =  n07 & ~n11;
assign n29 = ~n27 &  n28;
assign n30 = ~n26 &  n29;
assign n31 = ~n06 & ~n07;
assign n32 = ~n09 &  n31;
assign n33 = ~n05 &  n08;
assign n34 = ~n10 & ~n33;
assign n35 = ~n32 & ~n34;
assign n36 = ~n30 &  n35;
assign n37 = ~n12 & ~n36;
assign n38 =  n01 &  n03;
assign n39 = ~n11 &  n19;
assign n40 = ~n05 & ~n06;
assign n41 = ~n39 &  n40;
assign n42 = ~n38 & ~n41;
assign n43 =  n08 & ~n11;
assign n44 =  n05 & ~n12;
assign n45 = ~n43 & ~n44;
assign n46 =  n31 & ~n45;
assign n47 =  n01 &  n04;
assign n48 =  n02 &  n03;
assign n49 =  n07 & ~n48;
assign n50 = ~n47 &  n49;
assign n51 = ~n46 & ~n50;
assign n52 = ~n42 &  n51;
assign n53 = ~n37 &  n52;
assign n54 = ~n25 &  n53;
assign n17 =  n54;
endmodule

